library verilog;
use verilog.vl_types.all;
entity testbench_timer is
end testbench_timer;
